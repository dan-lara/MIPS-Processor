module alu (
	input 	  [31:0] EntradaA, EntradaB,
	input 	  [1:0] OP,
	output reg [31:0] Saida
);

	always @(*)begin
		case(OP)
			2'b00: Saida <= EntradaA + EntradaB;
			2'b01: Saida <= EntradaA - EntradaB;
			2'b10: Saida <= EntradaA & EntradaB;
			2'b11: Saida <= EntradaA | EntradaB;
		endcase
	end
endmodule	